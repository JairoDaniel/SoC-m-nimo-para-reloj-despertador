// taller.v

// Generated using ACDS version 18.0 614

`timescale 1 ps / 1 ps
module taller (
		input  wire       button1_export, // button1.export
		input  wire       button2_export, // button2.export
		input  wire       button3_export, // button3.export
		input  wire       clk_clk,        //     clk.clk
		output wire [7:0] leds_export,    //    leds.export
		input  wire       reset_reset_n,  //   reset.reset_n
		output wire [6:0] seg1_export,    //    seg1.export
		output wire [6:0] seg2_export,    //    seg2.export
		output wire [6:0] seg3_export,    //    seg3.export
		output wire [6:0] seg4_export,    //    seg4.export
		input  wire       uart_rxd,       //    uart.rxd
		output wire       uart_txd        //        .txd
	);

	wire  [31:0] cpu_data_master_readdata;                             // mm_interconnect_0:CPU_data_master_readdata -> CPU:d_readdata
	wire         cpu_data_master_waitrequest;                          // mm_interconnect_0:CPU_data_master_waitrequest -> CPU:d_waitrequest
	wire         cpu_data_master_debugaccess;                          // CPU:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:CPU_data_master_debugaccess
	wire  [15:0] cpu_data_master_address;                              // CPU:d_address -> mm_interconnect_0:CPU_data_master_address
	wire   [3:0] cpu_data_master_byteenable;                           // CPU:d_byteenable -> mm_interconnect_0:CPU_data_master_byteenable
	wire         cpu_data_master_read;                                 // CPU:d_read -> mm_interconnect_0:CPU_data_master_read
	wire         cpu_data_master_write;                                // CPU:d_write -> mm_interconnect_0:CPU_data_master_write
	wire  [31:0] cpu_data_master_writedata;                            // CPU:d_writedata -> mm_interconnect_0:CPU_data_master_writedata
	wire  [31:0] cpu_instruction_master_readdata;                      // mm_interconnect_0:CPU_instruction_master_readdata -> CPU:i_readdata
	wire         cpu_instruction_master_waitrequest;                   // mm_interconnect_0:CPU_instruction_master_waitrequest -> CPU:i_waitrequest
	wire  [15:0] cpu_instruction_master_address;                       // CPU:i_address -> mm_interconnect_0:CPU_instruction_master_address
	wire         cpu_instruction_master_read;                          // CPU:i_read -> mm_interconnect_0:CPU_instruction_master_read
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;  // mm_interconnect_0:JTAG_avalon_jtag_slave_chipselect -> JTAG:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;    // JTAG:av_readdata -> mm_interconnect_0:JTAG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest; // JTAG:av_waitrequest -> mm_interconnect_0:JTAG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;     // mm_interconnect_0:JTAG_avalon_jtag_slave_address -> JTAG:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;        // mm_interconnect_0:JTAG_avalon_jtag_slave_read -> JTAG:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;       // mm_interconnect_0:JTAG_avalon_jtag_slave_write -> JTAG:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;   // mm_interconnect_0:JTAG_avalon_jtag_slave_writedata -> JTAG:av_writedata
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_readdata;       // CPU:debug_mem_slave_readdata -> mm_interconnect_0:CPU_debug_mem_slave_readdata
	wire         mm_interconnect_0_cpu_debug_mem_slave_waitrequest;    // CPU:debug_mem_slave_waitrequest -> mm_interconnect_0:CPU_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_cpu_debug_mem_slave_debugaccess;    // mm_interconnect_0:CPU_debug_mem_slave_debugaccess -> CPU:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_cpu_debug_mem_slave_address;        // mm_interconnect_0:CPU_debug_mem_slave_address -> CPU:debug_mem_slave_address
	wire         mm_interconnect_0_cpu_debug_mem_slave_read;           // mm_interconnect_0:CPU_debug_mem_slave_read -> CPU:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_cpu_debug_mem_slave_byteenable;     // mm_interconnect_0:CPU_debug_mem_slave_byteenable -> CPU:debug_mem_slave_byteenable
	wire         mm_interconnect_0_cpu_debug_mem_slave_write;          // mm_interconnect_0:CPU_debug_mem_slave_write -> CPU:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_cpu_debug_mem_slave_writedata;      // mm_interconnect_0:CPU_debug_mem_slave_writedata -> CPU:debug_mem_slave_writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                  // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                    // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [11:0] mm_interconnect_0_ram_s1_address;                     // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                  // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                       // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                   // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                       // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         mm_interconnect_0_leds_s1_chipselect;                 // mm_interconnect_0:LEDS_s1_chipselect -> LEDS:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                   // LEDS:readdata -> mm_interconnect_0:LEDS_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                    // mm_interconnect_0:LEDS_s1_address -> LEDS:address
	wire         mm_interconnect_0_leds_s1_write;                      // mm_interconnect_0:LEDS_s1_write -> LEDS:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                  // mm_interconnect_0:LEDS_s1_writedata -> LEDS:writedata
	wire         mm_interconnect_0_seg1_s1_chipselect;                 // mm_interconnect_0:SEG1_s1_chipselect -> SEG1:chipselect
	wire  [31:0] mm_interconnect_0_seg1_s1_readdata;                   // SEG1:readdata -> mm_interconnect_0:SEG1_s1_readdata
	wire   [2:0] mm_interconnect_0_seg1_s1_address;                    // mm_interconnect_0:SEG1_s1_address -> SEG1:address
	wire         mm_interconnect_0_seg1_s1_write;                      // mm_interconnect_0:SEG1_s1_write -> SEG1:write_n
	wire  [31:0] mm_interconnect_0_seg1_s1_writedata;                  // mm_interconnect_0:SEG1_s1_writedata -> SEG1:writedata
	wire         mm_interconnect_0_button1_s1_chipselect;              // mm_interconnect_0:BUTTON1_s1_chipselect -> BUTTON1:chipselect
	wire  [31:0] mm_interconnect_0_button1_s1_readdata;                // BUTTON1:readdata -> mm_interconnect_0:BUTTON1_s1_readdata
	wire   [1:0] mm_interconnect_0_button1_s1_address;                 // mm_interconnect_0:BUTTON1_s1_address -> BUTTON1:address
	wire         mm_interconnect_0_button1_s1_write;                   // mm_interconnect_0:BUTTON1_s1_write -> BUTTON1:write_n
	wire  [31:0] mm_interconnect_0_button1_s1_writedata;               // mm_interconnect_0:BUTTON1_s1_writedata -> BUTTON1:writedata
	wire         mm_interconnect_0_timer_s1_chipselect;                // mm_interconnect_0:TIMER_s1_chipselect -> TIMER:chipselect
	wire  [15:0] mm_interconnect_0_timer_s1_readdata;                  // TIMER:readdata -> mm_interconnect_0:TIMER_s1_readdata
	wire   [2:0] mm_interconnect_0_timer_s1_address;                   // mm_interconnect_0:TIMER_s1_address -> TIMER:address
	wire         mm_interconnect_0_timer_s1_write;                     // mm_interconnect_0:TIMER_s1_write -> TIMER:write_n
	wire  [15:0] mm_interconnect_0_timer_s1_writedata;                 // mm_interconnect_0:TIMER_s1_writedata -> TIMER:writedata
	wire         mm_interconnect_0_button2_s1_chipselect;              // mm_interconnect_0:BUTTON2_s1_chipselect -> BUTTON2:chipselect
	wire  [31:0] mm_interconnect_0_button2_s1_readdata;                // BUTTON2:readdata -> mm_interconnect_0:BUTTON2_s1_readdata
	wire   [1:0] mm_interconnect_0_button2_s1_address;                 // mm_interconnect_0:BUTTON2_s1_address -> BUTTON2:address
	wire         mm_interconnect_0_button2_s1_write;                   // mm_interconnect_0:BUTTON2_s1_write -> BUTTON2:write_n
	wire  [31:0] mm_interconnect_0_button2_s1_writedata;               // mm_interconnect_0:BUTTON2_s1_writedata -> BUTTON2:writedata
	wire         mm_interconnect_0_button3_s1_chipselect;              // mm_interconnect_0:BUTTON3_s1_chipselect -> BUTTON3:chipselect
	wire  [31:0] mm_interconnect_0_button3_s1_readdata;                // BUTTON3:readdata -> mm_interconnect_0:BUTTON3_s1_readdata
	wire   [1:0] mm_interconnect_0_button3_s1_address;                 // mm_interconnect_0:BUTTON3_s1_address -> BUTTON3:address
	wire         mm_interconnect_0_button3_s1_write;                   // mm_interconnect_0:BUTTON3_s1_write -> BUTTON3:write_n
	wire  [31:0] mm_interconnect_0_button3_s1_writedata;               // mm_interconnect_0:BUTTON3_s1_writedata -> BUTTON3:writedata
	wire         mm_interconnect_0_seg2_s1_chipselect;                 // mm_interconnect_0:SEG2_s1_chipselect -> SEG2:chipselect
	wire  [31:0] mm_interconnect_0_seg2_s1_readdata;                   // SEG2:readdata -> mm_interconnect_0:SEG2_s1_readdata
	wire   [1:0] mm_interconnect_0_seg2_s1_address;                    // mm_interconnect_0:SEG2_s1_address -> SEG2:address
	wire         mm_interconnect_0_seg2_s1_write;                      // mm_interconnect_0:SEG2_s1_write -> SEG2:write_n
	wire  [31:0] mm_interconnect_0_seg2_s1_writedata;                  // mm_interconnect_0:SEG2_s1_writedata -> SEG2:writedata
	wire         mm_interconnect_0_seg3_s1_chipselect;                 // mm_interconnect_0:SEG3_s1_chipselect -> SEG3:chipselect
	wire  [31:0] mm_interconnect_0_seg3_s1_readdata;                   // SEG3:readdata -> mm_interconnect_0:SEG3_s1_readdata
	wire   [1:0] mm_interconnect_0_seg3_s1_address;                    // mm_interconnect_0:SEG3_s1_address -> SEG3:address
	wire         mm_interconnect_0_seg3_s1_write;                      // mm_interconnect_0:SEG3_s1_write -> SEG3:write_n
	wire  [31:0] mm_interconnect_0_seg3_s1_writedata;                  // mm_interconnect_0:SEG3_s1_writedata -> SEG3:writedata
	wire         mm_interconnect_0_seg4_s1_chipselect;                 // mm_interconnect_0:SEG4_s1_chipselect -> SEG4:chipselect
	wire  [31:0] mm_interconnect_0_seg4_s1_readdata;                   // SEG4:readdata -> mm_interconnect_0:SEG4_s1_readdata
	wire   [1:0] mm_interconnect_0_seg4_s1_address;                    // mm_interconnect_0:SEG4_s1_address -> SEG4:address
	wire         mm_interconnect_0_seg4_s1_write;                      // mm_interconnect_0:SEG4_s1_write -> SEG4:write_n
	wire  [31:0] mm_interconnect_0_seg4_s1_writedata;                  // mm_interconnect_0:SEG4_s1_writedata -> SEG4:writedata
	wire         mm_interconnect_0_uart_s1_chipselect;                 // mm_interconnect_0:UART_s1_chipselect -> UART:chipselect
	wire  [15:0] mm_interconnect_0_uart_s1_readdata;                   // UART:readdata -> mm_interconnect_0:UART_s1_readdata
	wire   [2:0] mm_interconnect_0_uart_s1_address;                    // mm_interconnect_0:UART_s1_address -> UART:address
	wire         mm_interconnect_0_uart_s1_read;                       // mm_interconnect_0:UART_s1_read -> UART:read_n
	wire         mm_interconnect_0_uart_s1_begintransfer;              // mm_interconnect_0:UART_s1_begintransfer -> UART:begintransfer
	wire         mm_interconnect_0_uart_s1_write;                      // mm_interconnect_0:UART_s1_write -> UART:write_n
	wire  [15:0] mm_interconnect_0_uart_s1_writedata;                  // mm_interconnect_0:UART_s1_writedata -> UART:writedata
	wire         irq_mapper_receiver0_irq;                             // JTAG:av_irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                             // BUTTON1:irq -> irq_mapper:receiver1_irq
	wire         irq_mapper_receiver2_irq;                             // TIMER:irq -> irq_mapper:receiver2_irq
	wire         irq_mapper_receiver3_irq;                             // BUTTON2:irq -> irq_mapper:receiver3_irq
	wire         irq_mapper_receiver4_irq;                             // BUTTON3:irq -> irq_mapper:receiver4_irq
	wire         irq_mapper_receiver5_irq;                             // UART:irq -> irq_mapper:receiver5_irq
	wire  [31:0] cpu_irq_irq;                                          // irq_mapper:sender_irq -> CPU:irq
	wire         rst_controller_reset_out_reset;                       // rst_controller:reset_out -> [BUTTON1:reset_n, BUTTON2:reset_n, BUTTON3:reset_n, UART:reset_n, mm_interconnect_0:BUTTON1_reset_reset_bridge_in_reset_reset]
	wire         cpu_debug_reset_request_reset;                        // CPU:debug_reset_request -> rst_controller:reset_in1
	wire         rst_controller_001_reset_out_reset;                   // rst_controller_001:reset_out -> [CPU:reset_n, JTAG:rst_n, LEDS:reset_n, RAM:reset, SEG1:reset_n, SEG2:reset_n, SEG3:reset_n, SEG4:reset_n, TIMER:reset_n, irq_mapper:reset, mm_interconnect_0:CPU_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_001_reset_out_reset_req;               // rst_controller_001:reset_req -> [CPU:reset_req, RAM:reset_req, rst_translator:reset_req_in]

	taller_BUTTON1 button1 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_button1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button1_s1_readdata),   //                    .readdata
		.in_port    (button1_export),                          // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                 //                 irq.irq
	);

	taller_BUTTON1 button2 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_button2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button2_s1_readdata),   //                    .readdata
		.in_port    (button2_export),                          // external_connection.export
		.irq        (irq_mapper_receiver3_irq)                 //                 irq.irq
	);

	taller_BUTTON1 button3 (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_button3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_button3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_button3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_button3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_button3_s1_readdata),   //                    .readdata
		.in_port    (button3_export),                          // external_connection.export
		.irq        (irq_mapper_receiver4_irq)                 //                 irq.irq
	);

	taller_CPU cpu (
		.clk                                 (clk_clk),                                           //                       clk.clk
		.reset_n                             (~rst_controller_001_reset_out_reset),               //                     reset.reset_n
		.reset_req                           (rst_controller_001_reset_out_reset_req),            //                          .reset_req
		.d_address                           (cpu_data_master_address),                           //               data_master.address
		.d_byteenable                        (cpu_data_master_byteenable),                        //                          .byteenable
		.d_read                              (cpu_data_master_read),                              //                          .read
		.d_readdata                          (cpu_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (cpu_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (cpu_data_master_write),                             //                          .write
		.d_writedata                         (cpu_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (cpu_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (cpu_instruction_master_address),                    //        instruction_master.address
		.i_read                              (cpu_instruction_master_read),                       //                          .read
		.i_readdata                          (cpu_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (cpu_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (cpu_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (cpu_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_cpu_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_cpu_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_cpu_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_cpu_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_cpu_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_cpu_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_cpu_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_cpu_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                   // custom_instruction_master.readra
	);

	taller_JTAG jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_001_reset_out_reset),                  //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                              //               irq.irq
	);

	taller_LEDS leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	taller_RAM ram (
		.clk        (clk_clk),                                //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),       //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),         //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect),    //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),         //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),      //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),     //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable),    //       .byteenable
		.reset      (rst_controller_001_reset_out_reset),     // reset1.reset
		.reset_req  (rst_controller_001_reset_out_reset_req), //       .reset_req
		.freeze     (1'b0)                                    // (terminated)
	);

	taller_SEG1 seg1 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_0_seg1_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg1_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg1_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg1_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg1_s1_readdata),   //                    .readdata
		.out_port   (seg1_export)                           // external_connection.export
	);

	taller_SEG2 seg2 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_0_seg2_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg2_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg2_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg2_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg2_s1_readdata),   //                    .readdata
		.out_port   (seg2_export)                           // external_connection.export
	);

	taller_SEG2 seg3 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_0_seg3_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg3_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg3_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg3_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg3_s1_readdata),   //                    .readdata
		.out_port   (seg3_export)                           // external_connection.export
	);

	taller_SEG2 seg4 (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_001_reset_out_reset),  //               reset.reset_n
		.address    (mm_interconnect_0_seg4_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_seg4_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_seg4_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_seg4_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_seg4_s1_readdata),   //                    .readdata
		.out_port   (seg4_export)                           // external_connection.export
	);

	taller_TIMER timer (
		.clk           (clk_clk),                               //           clk.clk
		.reset_n       (~rst_controller_001_reset_out_reset),   //         reset.reset_n
		.address       (mm_interconnect_0_timer_s1_address),    //            s1.address
		.writedata     (mm_interconnect_0_timer_s1_writedata),  //              .writedata
		.readdata      (mm_interconnect_0_timer_s1_readdata),   //              .readdata
		.chipselect    (mm_interconnect_0_timer_s1_chipselect), //              .chipselect
		.write_n       (~mm_interconnect_0_timer_s1_write),     //              .write_n
		.irq           (irq_mapper_receiver2_irq),              //           irq.irq
		.timeout_pulse ()                                       // external_port.export
	);

	taller_UART uart (
		.clk           (clk_clk),                                 //                 clk.clk
		.reset_n       (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address       (mm_interconnect_0_uart_s1_address),       //                  s1.address
		.begintransfer (mm_interconnect_0_uart_s1_begintransfer), //                    .begintransfer
		.chipselect    (mm_interconnect_0_uart_s1_chipselect),    //                    .chipselect
		.read_n        (~mm_interconnect_0_uart_s1_read),         //                    .read_n
		.write_n       (~mm_interconnect_0_uart_s1_write),        //                    .write_n
		.writedata     (mm_interconnect_0_uart_s1_writedata),     //                    .writedata
		.readdata      (mm_interconnect_0_uart_s1_readdata),      //                    .readdata
		.rxd           (uart_rxd),                                // external_connection.export
		.txd           (uart_txd),                                //                    .export
		.irq           (irq_mapper_receiver5_irq)                 //                 irq.irq
	);

	taller_mm_interconnect_0 mm_interconnect_0 (
		.CLOCK_clk_clk                             (clk_clk),                                              //                           CLOCK_clk.clk
		.BUTTON1_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                       // BUTTON1_reset_reset_bridge_in_reset.reset
		.CPU_reset_reset_bridge_in_reset_reset     (rst_controller_001_reset_out_reset),                   //     CPU_reset_reset_bridge_in_reset.reset
		.CPU_data_master_address                   (cpu_data_master_address),                              //                     CPU_data_master.address
		.CPU_data_master_waitrequest               (cpu_data_master_waitrequest),                          //                                    .waitrequest
		.CPU_data_master_byteenable                (cpu_data_master_byteenable),                           //                                    .byteenable
		.CPU_data_master_read                      (cpu_data_master_read),                                 //                                    .read
		.CPU_data_master_readdata                  (cpu_data_master_readdata),                             //                                    .readdata
		.CPU_data_master_write                     (cpu_data_master_write),                                //                                    .write
		.CPU_data_master_writedata                 (cpu_data_master_writedata),                            //                                    .writedata
		.CPU_data_master_debugaccess               (cpu_data_master_debugaccess),                          //                                    .debugaccess
		.CPU_instruction_master_address            (cpu_instruction_master_address),                       //              CPU_instruction_master.address
		.CPU_instruction_master_waitrequest        (cpu_instruction_master_waitrequest),                   //                                    .waitrequest
		.CPU_instruction_master_read               (cpu_instruction_master_read),                          //                                    .read
		.CPU_instruction_master_readdata           (cpu_instruction_master_readdata),                      //                                    .readdata
		.BUTTON1_s1_address                        (mm_interconnect_0_button1_s1_address),                 //                          BUTTON1_s1.address
		.BUTTON1_s1_write                          (mm_interconnect_0_button1_s1_write),                   //                                    .write
		.BUTTON1_s1_readdata                       (mm_interconnect_0_button1_s1_readdata),                //                                    .readdata
		.BUTTON1_s1_writedata                      (mm_interconnect_0_button1_s1_writedata),               //                                    .writedata
		.BUTTON1_s1_chipselect                     (mm_interconnect_0_button1_s1_chipselect),              //                                    .chipselect
		.BUTTON2_s1_address                        (mm_interconnect_0_button2_s1_address),                 //                          BUTTON2_s1.address
		.BUTTON2_s1_write                          (mm_interconnect_0_button2_s1_write),                   //                                    .write
		.BUTTON2_s1_readdata                       (mm_interconnect_0_button2_s1_readdata),                //                                    .readdata
		.BUTTON2_s1_writedata                      (mm_interconnect_0_button2_s1_writedata),               //                                    .writedata
		.BUTTON2_s1_chipselect                     (mm_interconnect_0_button2_s1_chipselect),              //                                    .chipselect
		.BUTTON3_s1_address                        (mm_interconnect_0_button3_s1_address),                 //                          BUTTON3_s1.address
		.BUTTON3_s1_write                          (mm_interconnect_0_button3_s1_write),                   //                                    .write
		.BUTTON3_s1_readdata                       (mm_interconnect_0_button3_s1_readdata),                //                                    .readdata
		.BUTTON3_s1_writedata                      (mm_interconnect_0_button3_s1_writedata),               //                                    .writedata
		.BUTTON3_s1_chipselect                     (mm_interconnect_0_button3_s1_chipselect),              //                                    .chipselect
		.CPU_debug_mem_slave_address               (mm_interconnect_0_cpu_debug_mem_slave_address),        //                 CPU_debug_mem_slave.address
		.CPU_debug_mem_slave_write                 (mm_interconnect_0_cpu_debug_mem_slave_write),          //                                    .write
		.CPU_debug_mem_slave_read                  (mm_interconnect_0_cpu_debug_mem_slave_read),           //                                    .read
		.CPU_debug_mem_slave_readdata              (mm_interconnect_0_cpu_debug_mem_slave_readdata),       //                                    .readdata
		.CPU_debug_mem_slave_writedata             (mm_interconnect_0_cpu_debug_mem_slave_writedata),      //                                    .writedata
		.CPU_debug_mem_slave_byteenable            (mm_interconnect_0_cpu_debug_mem_slave_byteenable),     //                                    .byteenable
		.CPU_debug_mem_slave_waitrequest           (mm_interconnect_0_cpu_debug_mem_slave_waitrequest),    //                                    .waitrequest
		.CPU_debug_mem_slave_debugaccess           (mm_interconnect_0_cpu_debug_mem_slave_debugaccess),    //                                    .debugaccess
		.JTAG_avalon_jtag_slave_address            (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //              JTAG_avalon_jtag_slave.address
		.JTAG_avalon_jtag_slave_write              (mm_interconnect_0_jtag_avalon_jtag_slave_write),       //                                    .write
		.JTAG_avalon_jtag_slave_read               (mm_interconnect_0_jtag_avalon_jtag_slave_read),        //                                    .read
		.JTAG_avalon_jtag_slave_readdata           (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                                    .readdata
		.JTAG_avalon_jtag_slave_writedata          (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                                    .writedata
		.JTAG_avalon_jtag_slave_waitrequest        (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                                    .waitrequest
		.JTAG_avalon_jtag_slave_chipselect         (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  //                                    .chipselect
		.LEDS_s1_address                           (mm_interconnect_0_leds_s1_address),                    //                             LEDS_s1.address
		.LEDS_s1_write                             (mm_interconnect_0_leds_s1_write),                      //                                    .write
		.LEDS_s1_readdata                          (mm_interconnect_0_leds_s1_readdata),                   //                                    .readdata
		.LEDS_s1_writedata                         (mm_interconnect_0_leds_s1_writedata),                  //                                    .writedata
		.LEDS_s1_chipselect                        (mm_interconnect_0_leds_s1_chipselect),                 //                                    .chipselect
		.RAM_s1_address                            (mm_interconnect_0_ram_s1_address),                     //                              RAM_s1.address
		.RAM_s1_write                              (mm_interconnect_0_ram_s1_write),                       //                                    .write
		.RAM_s1_readdata                           (mm_interconnect_0_ram_s1_readdata),                    //                                    .readdata
		.RAM_s1_writedata                          (mm_interconnect_0_ram_s1_writedata),                   //                                    .writedata
		.RAM_s1_byteenable                         (mm_interconnect_0_ram_s1_byteenable),                  //                                    .byteenable
		.RAM_s1_chipselect                         (mm_interconnect_0_ram_s1_chipselect),                  //                                    .chipselect
		.RAM_s1_clken                              (mm_interconnect_0_ram_s1_clken),                       //                                    .clken
		.SEG1_s1_address                           (mm_interconnect_0_seg1_s1_address),                    //                             SEG1_s1.address
		.SEG1_s1_write                             (mm_interconnect_0_seg1_s1_write),                      //                                    .write
		.SEG1_s1_readdata                          (mm_interconnect_0_seg1_s1_readdata),                   //                                    .readdata
		.SEG1_s1_writedata                         (mm_interconnect_0_seg1_s1_writedata),                  //                                    .writedata
		.SEG1_s1_chipselect                        (mm_interconnect_0_seg1_s1_chipselect),                 //                                    .chipselect
		.SEG2_s1_address                           (mm_interconnect_0_seg2_s1_address),                    //                             SEG2_s1.address
		.SEG2_s1_write                             (mm_interconnect_0_seg2_s1_write),                      //                                    .write
		.SEG2_s1_readdata                          (mm_interconnect_0_seg2_s1_readdata),                   //                                    .readdata
		.SEG2_s1_writedata                         (mm_interconnect_0_seg2_s1_writedata),                  //                                    .writedata
		.SEG2_s1_chipselect                        (mm_interconnect_0_seg2_s1_chipselect),                 //                                    .chipselect
		.SEG3_s1_address                           (mm_interconnect_0_seg3_s1_address),                    //                             SEG3_s1.address
		.SEG3_s1_write                             (mm_interconnect_0_seg3_s1_write),                      //                                    .write
		.SEG3_s1_readdata                          (mm_interconnect_0_seg3_s1_readdata),                   //                                    .readdata
		.SEG3_s1_writedata                         (mm_interconnect_0_seg3_s1_writedata),                  //                                    .writedata
		.SEG3_s1_chipselect                        (mm_interconnect_0_seg3_s1_chipselect),                 //                                    .chipselect
		.SEG4_s1_address                           (mm_interconnect_0_seg4_s1_address),                    //                             SEG4_s1.address
		.SEG4_s1_write                             (mm_interconnect_0_seg4_s1_write),                      //                                    .write
		.SEG4_s1_readdata                          (mm_interconnect_0_seg4_s1_readdata),                   //                                    .readdata
		.SEG4_s1_writedata                         (mm_interconnect_0_seg4_s1_writedata),                  //                                    .writedata
		.SEG4_s1_chipselect                        (mm_interconnect_0_seg4_s1_chipselect),                 //                                    .chipselect
		.TIMER_s1_address                          (mm_interconnect_0_timer_s1_address),                   //                            TIMER_s1.address
		.TIMER_s1_write                            (mm_interconnect_0_timer_s1_write),                     //                                    .write
		.TIMER_s1_readdata                         (mm_interconnect_0_timer_s1_readdata),                  //                                    .readdata
		.TIMER_s1_writedata                        (mm_interconnect_0_timer_s1_writedata),                 //                                    .writedata
		.TIMER_s1_chipselect                       (mm_interconnect_0_timer_s1_chipselect),                //                                    .chipselect
		.UART_s1_address                           (mm_interconnect_0_uart_s1_address),                    //                             UART_s1.address
		.UART_s1_write                             (mm_interconnect_0_uart_s1_write),                      //                                    .write
		.UART_s1_read                              (mm_interconnect_0_uart_s1_read),                       //                                    .read
		.UART_s1_readdata                          (mm_interconnect_0_uart_s1_readdata),                   //                                    .readdata
		.UART_s1_writedata                         (mm_interconnect_0_uart_s1_writedata),                  //                                    .writedata
		.UART_s1_begintransfer                     (mm_interconnect_0_uart_s1_begintransfer),              //                                    .begintransfer
		.UART_s1_chipselect                        (mm_interconnect_0_uart_s1_chipselect)                  //                                    .chipselect
	);

	taller_irq_mapper irq_mapper (
		.clk           (clk_clk),                            //       clk.clk
		.reset         (rst_controller_001_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.receiver5_irq (irq_mapper_receiver5_irq),           // receiver5.irq
		.sender_irq    (cpu_irq_irq)                         //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.reset_in1      (cpu_debug_reset_request_reset),  // reset_in1.reset
		.clk            (clk_clk),                        //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                         // reset_in0.reset
		.clk            (clk_clk),                                //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_001_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_in1      (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

endmodule
